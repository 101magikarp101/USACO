// TODO: Implement the basic pipeline module
// This module should implement a 5-stage pipeline for arithmetic operations
// Stages: Fetch, Decode, Execute, Memory, Writeback
// The pipeline should take two 8-bit inputs and produce an 8-bit result

module pipeline_arith (
  input         clk,
  input         rst,
  input  [7:0]  a,
  input  [7:0]  b,
  output reg [7:0] result
);
  // Your implementation here
  
endmodule
